LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULTIPLIER32_toplevel IS
   PORT (--

        inA               : IN std_logic_vector(31 DOWNTO 0);
        inB               : IN std_logic_vector(31 DOWNTO 0);
	start		  : IN std_logic;
	clk		  : IN std_logic;
	clear		  : IN std_logic;

	output		  : OUT std_logic_vector(63 DOWNTO 0);
	done		  : OUT std_logic
   );
END MULTIPLIER32_toplevel;

ARCHITECTURE struct OF MULTIPLIER32_toplevel IS



--MULTIPLIER32_toplevel has a 5 bit counter, 3 32 bit shift register, 2 flip-flops, 32 bit adder, 32bit xor, MUL32_controller

COMPONENT XOR32 IS
   PORT (--

        in32               : IN std_logic_vector(31 DOWNTO 0);
	control2s	  : IN std_logic; -- control2s=1, 1's compliment, or what it is
        Out32               : OUT std_logic_vector(31 DOWNTO 0)

   );
END COMPONENT;

COMPONENT COUNTER_5BIT IS
   PORT (--
         clk                : IN std_logic;
         en                : IN std_logic;
	 clear             : IN std_logic; 

         q                : OUT std_logic_vector(4 DOWNTO 0);
	 over		  : OUT std_logic

   );
END COMPONENT;

COMPONENT SHIFT_32bit IS
   PORT (--
	hold		  : IN std_logic;
        sin               : IN std_logic;
        pin               : IN std_logic_vector(31 DOWNTO 0);
	ld_shiftb	  : IN std_logic;
	clk		  : IN std_logic;
	clear		  : IN std_logic;
	qsout 		  : OUT std_logic; --serial out
	qpout		  : OUT std_logic_vector(31 DOWNTO 0)
   );
END COMPONENT;

COMPONENT DFF_DTFL IS
   PORT (--
         d                : IN std_logic;
         clk                : IN std_logic;
	 clear			: IN std_logic;	

	 q 		    : OUT std_logic
   );
END COMPONENT;

COMPONENT FULLADDER33bit IS
   PORT (--
         
	x	: IN std_logic_vector(32 DOWNTO 0);    
	y	: IN std_logic_vector(32 DOWNTO 0);
	cin	: IN std_logic;         
	sum     : OUT std_logic_vector(32 DOWNTO 0);
	cout    : OUT std_logic
   );
END COMPONENT;

COMPONENT MUL32_controller IS
   PORT(
	start		   : IN std_logic;
	a		   : IN std_logic_vector(1 DOWNTO 0);
	cnt_done	   : IN std_logic;
	clk		   : IN std_logic;
	clear		   : IN std_logic;

	done		   : OUT std_logic;
	control2s	   : OUT std_logic;
	hold32		   : OUT std_logic;
	hold33		   : OUT std_logic;
	holdX		   : OUT std_logic;
	ld_rshiftb	   : OUT std_logic;
	counter_en	   : OUT std_logic;
	counter_clear	   : OUT std_logic;
	muxout		   : OUT std_logic);
END COMPONENT;




COMPONENT MUX33bit1sel IS
   PORT (--
         in0                : IN std_logic_vector(32 DOWNTO 0);
         in1                : IN std_logic_vector(32 DOWNTO 0);
	
         s0                : IN std_logic;

	 out33 		    : OUT std_logic_vector(32 DOWNTO 0)
   );
END COMPONENT;

COMPONENT SHIFT_33bit IS
   PORT (--
	hold		  : IN std_logic;
        sin               : IN std_logic;
        pin               : IN std_logic_vector(32 DOWNTO 0);
	ld_shiftb	  : IN std_logic;
	clk		  : IN std_logic;
	clear		  : IN std_logic;
	qsout 		  : OUT std_logic; --serial out
	qpout		  : OUT std_logic_vector(32 DOWNTO 0)
   );
END COMPONENT;

COMPONENT MUX2to1 IS
   PORT (--
         in0                : IN std_logic;
         in1                : IN std_logic;
	
         s0                : IN std_logic;

	 out2to1 		    : OUT std_logic
   );
END COMPONENT;
--binding

FOR ALL: XOR32 USE ENTITY WORK.XOR32(struct);
FOR ALL: MUX2to1 USE ENTITY WORK.MUX2to1(struct);
FOR ALL: SHIFT_32bit USE ENTITY WORK.SHIFT_32bit(struct);
FOR ALL: MUL32_controller USE ENTITY WORK.MUL32_controller(behav);
FOR ALL: DFF_DTFL USE ENTITY WORK.DFF_DTFL(dataflow);
FOR ALL: FULLADDER33bit USE ENTITY WORK.FULLADDER33bit(struct);
FOR ALL: COUNTER_5BIT USE ENTITY WORK.COUNTER_5BIT(struct);
--FOR ALL: AND5 USE ENTITY WORK.AND5(dataflow);
FOR ALL: MUX33bit1sel USE ENTITY WORK.MUX33bit1sel(behav);

FOR ALL: SHIFT_33bit USE ENTITY WORK.SHIFT_33bit(struct);


--temp signal for the 4 branches
SIGNAL tempAllZeros : std_logic_vector(32 DOWNTO 0):="000000000000000000000000000000000";
SIGNAL tempP, tempB2, tempmAdder, tempXAdder, tempAdder: std_logic_vector(32 DOWNTO 0);--:="000000000000000000000000000000000";
SIGNAL tempA, tempB1 :std_logic_vector(31 DOWNTO 0);--:="00000000000000000000000000000000";
SIGNAL temps1, temps2, temps3, temps4, temps7, tempC	: std_logic:='0';
SIGNAL hold32, hold33, holdX, ld_shiftb, counter_en, counter_clear, control2s, done_t, cnt_done, start_t, muxout  : std_logic:='0';
SIGNAL tempZero: std_logic := '0';
SIGNAL tempOne: std_logic :='1';
SIGNAL temps5: std_logic:='0';
SIGNAL counter_out: std_logic_vector(4 DOWNTO 0):="00000";
SIGNAL a: std_logic_vector(1 DOWNTO 0):="00";
SIGNAL clkb, cnt_done_i: std_logic;
SIGNAL temps11: std_logic;

--start of process
BEGIN

	C10: clkb<= NOT clk;	

	T11: SHIFT_33bit PORT MAP (hold33, tempP(31), tempmAdder(32 DOWNTO 0), ld_shiftb, clk, clear, temps1, tempP(32 DOWNTO 0));

	
	--P0: SHIFT_32bit PORT MAP (hold, temps4, tempmAdder(31 DOWNTO 0), ld_shiftb, clk, clear, temps1, tempP(31 DOWNTO 0));
	--P1: tempP(32)<= temps4;

	Q0: SHIFT_32bit PORT MAP (hold32, temps1, inA, ld_shiftb, clk, clear, temps2, tempA);
	
	Q3: MUX2to1 PORT MAP (temps2, tempZero, muxout, temps11);

	Q1: DFF_DTFL PORT MAP (temps11, clk, clear, temps3);

	A0: FULLADDER33bit PORT MAP (tempP, tempB2, control2s, tempAdder, tempC);
	--A1: DFF_DTFL PORT MAP (tempmAdder(32), clk, clear, temps4);

	X10: SHIFT_33bit PORT MAP (holdX, tempZero, tempAdder, ld_shiftb, clkb, clear, temps7, tempXAdder);

	N0: SHIFT_32bit PORT MAP (tempZero, tempZero, inB, tempOne, clk, clear, temps5, tempB1);
	N1: XOR32 PORT MAP (tempB1, control2s, tempB2(31 DOWNTO 0));
	N2: tempB2(32)<=tempB2(31);	

	Z0: COUNTER_5BIT PORT MAP (clk, counter_en, counter_clear, counter_out, cnt_done_i);

	--Z10: AND5 PORT MAP(counter_out(4),counter_out(3),counter_out(2),counter_out(1),counter_out(0), cnt_done);
	Z10: cnt_done <= cnt_done_i;

	C0: a(1)<=temps2;
	C1: a(0)<=temps3; 
	C2: MUL32_controller PORT MAP(start, a, cnt_done, clk, clear, done, control2s, hold32, hold33, holdX, ld_shiftb, counter_en, counter_clear, muxout);	

	--M1: tempmAdder<=tempAdder;
	M0: MUX33bit1sel PORT MAP (tempXAdder, tempAllZeros, muxout, tempmAdder);

	O0: output(31 DOWNTO 0)<= tempA;
	O1: output(63 DOWNTO 32)<= tempP(31 DOWNTO 0);
END struct; 






